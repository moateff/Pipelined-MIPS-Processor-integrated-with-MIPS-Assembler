module imem #(parameter MEMFILE = "memfile.dat")(
	input  [5:0]  a,
	output [31:0] rd
);

	reg [31:0] RAM [63:0];

	initial begin
		$readmemh(MEMFILE, RAM, 0, 6);
	end

	assign rd = RAM[a]; // word aligned
	
endmodule

